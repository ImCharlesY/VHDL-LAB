 library ieee;                    
 use  ieee.std_logic_1164.all;     
 use  ieee.std_logic_unsigned.all; 
 
 entity ComunicateWithB20 is
 port(
	dq:buffer std_logic;
	sample:out std_logic_vector(7 downto 0)
 );
 end entity;
 
 architecture behavior of ComunicateWithB20 is
 ----------------------Signal Declaration-------------------
 
 ---------------------End Signal Declaration-----------------
 
 begin
 
 end behavior;